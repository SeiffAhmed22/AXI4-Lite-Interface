module axi4_lite_slave #(
    parameters
) (
    ports
);
    
endmodule