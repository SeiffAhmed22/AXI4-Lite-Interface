module axi4_lite_top #(
    parameters
) (
    ports
);
    
endmodule