module axi4_lite_master #(
    parameters
) (
    ports
);
    
endmodule